

module Test(
    input clk,
    input rst
);
   


endmodule
